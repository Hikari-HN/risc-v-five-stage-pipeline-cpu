`timescale 1ns / 1ps
//立即数扩展（0扩展或符号位扩展）
module Imm_gen(
    input  logic [31:0] inst_code,
    output logic [31:0] imm_out
);

    // add your immediate extension logic here.

endmodule
